/******************************************************************************* 
 * Module   : friscv_pipelined_top
 * Project  : FRiscV
 * Author   : Tom Szymkowiak
 * Mod. Date: 07-Feb-2021
 *******************************************************************************
 * Description:
 * ============
 * Top level for the 5-stage pipelined implementation of the FRiscV CPU
 ******************************************************************************/
module friscv_pipelined_top (

);

endmodule // friscv_pipelined_top