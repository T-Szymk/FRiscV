--****************************************************************************** 
-- Module   : friscv_pkg
-- Project  : FRiscV
-- Author   : Tom Szymkowiak
-- Mod. Date: 28-Dec-2021
--******************************************************************************
-- Description:
-- ============
-- VHDL package containing definitions and values that are used within the 
-- friscv project.
--******************************************************************************
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE friscv_pkg IS 
  
  	CONSTANT ARCH : INTEGER := 32;

END friscv_pkg;